`ifndef CFS_APB_SEQUENCE_RW_SV
 `define CFS_APB_SEQUENCE_RW_SV

class cfs_apb_sequence_rw extends cfs_apb_sequence_base;
  
  //public members that we allow inline randomization in test class
  rand cfs_apb_addr addr;
  rand cfs_apb_data wr_data;
  
  `uvm_object_utils(cfs_apb_sequence_rw)
  
  function new(string name = "");
    super.new(name);
  endfunction
  
  virtual task body();
    
    //such that we cannot access item directly from test class as there we want only addr and data to be accessible
    cfs_apb_item_drv item;
    
    //Read
    `uvm_do_with(item, {
      dir == CFS_APB_READ;
      //addr of the item we are randomizing = addr value in this class
      addr == local::addr;
    });
    
    //Write
    `uvm_do_with(item, {
      dir == CFS_APB_WRITE;
      //addr of the item we are randomizing = addr value in this class
      addr == local::addr;
      data == wr_data;
    });
   
  endtask
  
endclass


`endif
